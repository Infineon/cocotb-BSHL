// **************************************************************************
//
//  Author      : See AUTHORS
//  Project     : cocotb-BSHL
//  COPYRIGHT (c) 2023-24, Infineon Technologies AG. All rights reserved.
//
//  *****************************************************************************

package my_uvm_pkg;

        import uvm_pkg::*;
        `include "uvm_macros.svh"
        `include "my_transaction.svh"
        `include "my_scoreboard.svh"
        `include "my_monitor.svh"
        `include "my_driver.svh"
        `include "my_sequencer.svh"
        `include "my_sequence.svh"
        `include "my_agent.svh"
        `include "my_env.svh"

endpackage : my_uvm_pkg

